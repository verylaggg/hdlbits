module top_module_p114 ();
endmodule
