module top_module_p41 ();
endmodule
