module top_module_p37 ();
endmodule
