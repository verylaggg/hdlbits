module top_module_p48 ();
endmodule
