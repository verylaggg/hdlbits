module top_module_p121 ();
endmodule
