module top_module_p108 ();
endmodule
