module top_module_p66 ();
endmodule
