module top_module_p45 ();
endmodule
