module top_module_p142 ();
endmodule
