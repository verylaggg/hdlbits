module top_module_p139 ();
endmodule
