module top_module_p116 ();
endmodule
