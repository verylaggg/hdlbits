module top_module_p138 ();
endmodule
