module top_module_p20 ();
endmodule
