module top_module_p169 ();
endmodule
