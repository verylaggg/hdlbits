module top_module_p126 ();
endmodule
