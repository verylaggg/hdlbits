module top_module_p117 ();
endmodule
