module top_module_p182 ();
endmodule
