module top_module_p35 ();
endmodule
