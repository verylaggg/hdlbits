module top_module_p113 ();
endmodule
