module top_module_p70 ();
endmodule
