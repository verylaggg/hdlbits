module top_module_p147 ();
endmodule
