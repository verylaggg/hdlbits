module top_module_p21 ();
endmodule
