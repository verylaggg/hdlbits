module top_module_p71 ();
endmodule
