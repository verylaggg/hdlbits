module top_module_p153 ();
endmodule
