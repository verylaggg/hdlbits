module top_module_p17 ();
endmodule
