module top_module_p54 ( input x, input y, output z );
    assign z = ~(x ^ y);
endmodule
