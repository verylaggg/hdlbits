module top_module_p33 ();
endmodule
