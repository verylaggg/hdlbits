module top_module_p145 ();
endmodule
