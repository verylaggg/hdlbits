module top_module_p81 ();
endmodule
