module top_module_p90 ();
endmodule
