module top_module_p155 ();
endmodule
