module top_module_p118 ();
endmodule
