module top_module_p78 ();
endmodule
