module top_module_p88 ();
endmodule
