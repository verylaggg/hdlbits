module top_module_p173 ();
endmodule
