module top_module_p127 ();
endmodule
