module top_module_p38 ();
endmodule
