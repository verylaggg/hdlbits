module top_module_p30 ();
endmodule
