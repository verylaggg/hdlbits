module top_module_p73 ();
endmodule
