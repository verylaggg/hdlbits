module top_module_p89 ();
endmodule
