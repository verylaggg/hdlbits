module top_module_p3( input in, output out );
	assign out = in;
endmodule