module top_module_p32 ();
endmodule
