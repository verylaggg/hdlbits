module top_module_p85 ();
endmodule
