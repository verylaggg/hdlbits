module top_module_p179 ();
endmodule
