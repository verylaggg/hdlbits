module top_module_p172 ();
endmodule
