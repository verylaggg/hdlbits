module top_module_p8( 
    input a, 
    input b, 
    output out );
    
    assign out = ~(a ^ b);

endmodule
