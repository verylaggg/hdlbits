module top_module_p40 ();
endmodule
