module top_module_p151 ();
endmodule
