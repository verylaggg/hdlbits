module top_module_p158 ();
endmodule
