module top_module_p132 ();
endmodule
