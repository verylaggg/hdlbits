module top_module_p162 ();
endmodule
