module top_module_p39 ();
endmodule
