module top_module_p46 ();
endmodule
