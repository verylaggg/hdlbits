module top_module_p16 ();
endmodule
