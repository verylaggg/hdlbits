module top_module_p160 ();
endmodule
