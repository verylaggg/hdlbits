module top_module_p24 ();
endmodule
