module top_module_p76 ();
endmodule
