module top_module_p148 ();
endmodule
