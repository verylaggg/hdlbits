module top_module_p2(
    output zero
);// Module body starts after semicolon
	wire zero;
	assign zero = 1'b0;
endmodule
