module top_module_p143 ();
endmodule
