module top_module_p13 ();
endmodule
