module top_module_p86 ();
endmodule
