module top_module_p55 ();
endmodule
