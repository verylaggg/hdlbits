module top_module_p97 ();
endmodule
