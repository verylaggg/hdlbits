module top_module_p171 ();
endmodule
