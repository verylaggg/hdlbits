module top_module_p152 ();
endmodule
