module top_module_p31 ();
endmodule
