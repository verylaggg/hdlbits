module top_module_p180 ();
endmodule
