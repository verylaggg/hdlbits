module top_module_p65 ();
endmodule
