module top_module_p115 ();
endmodule
