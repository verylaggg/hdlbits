module top_module_p12 ();
endmodule
