module top_module_p83 ();
endmodule
