module top_module_p163 ();
endmodule
