module top_module_p64 ();
endmodule
