module top_module_p36 ();
endmodule
