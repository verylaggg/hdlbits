module top_module_p141 ();
endmodule
