module top_module_p170 ();
endmodule
