module top_module_p149 ();
endmodule
