module top_module_p5( input in, output out );
    assign out = ~in;
endmodule