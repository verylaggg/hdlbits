module top_module_p144 ();
endmodule
