module top_module_p164 ();
endmodule
