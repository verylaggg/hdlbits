module top_module_p92 ();
endmodule
