module top_module_p168 ();
endmodule
