module top_module_p146 ();
endmodule
