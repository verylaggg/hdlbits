module top_module_p122 ();
endmodule
