module top_module_p125 ();
endmodule
