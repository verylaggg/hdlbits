module top_module_p98 ();
endmodule
