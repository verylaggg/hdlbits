module top_module_p84 ();
endmodule
