module top_module_p14 ();
endmodule
