module top_module_p15 ();
endmodule
