module top_module_p53 ();
endmodule
