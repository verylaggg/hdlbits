module top_module_p43 ();
endmodule
