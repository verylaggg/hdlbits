module top_module_p50 ();
endmodule
