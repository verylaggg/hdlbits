module top_module_p77 ();
endmodule
