module top_module_p74 ();
endmodule
