module top_module_p1( output one );

// Insert your code here
    assign one = 1'b1;

endmodule