module top_module_p63 ();
endmodule
