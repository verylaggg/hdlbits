module top_module_p11 ();
endmodule
