module top_module_p112 ();
endmodule
