module top_module_p18 ();
endmodule
