module top_module_p93 ();
endmodule
