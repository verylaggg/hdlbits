module top_module_p6( 
    input a, 
    input b, 
    output out );
assign out = a & b;
endmodule