module top_module_p75 ();
endmodule
