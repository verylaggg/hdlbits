module top_module_p166 ();
endmodule
