module top_module_p23 ();
endmodule
