module top_module_p120 ();
endmodule
