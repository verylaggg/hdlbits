module top_module_p87 ();
endmodule
