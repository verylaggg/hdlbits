module top_module_p22 ();
endmodule
