module top_module_p150 ();
endmodule
