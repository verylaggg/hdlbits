module top_module_p52 ();
endmodule
