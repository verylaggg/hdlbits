module top_module_p140 ();
endmodule
