module top_module_p80 ();
endmodule
