//`define USE_DIY
module top_module ( 
    input [15:0] a, b,
    input cin,
    output cout,
    output [15:0] sum );
    wire [2:0]out;
`ifdef USE_DIY
    bcd_fadd_diy bcd_fadd0 (.a(a[3:0]), .b(b[3:0]), .cin(cin), .cout(out[0]), .sum(sum[3:0]));
    bcd_fadd_diy bcd_fadd1 (.a(a[7:4]), .b(b[7:4]), .cin(out[0]), .cout(out[1]), .sum(sum[7:4]));
    bcd_fadd_diy bcd_fadd2 (.a(a[11:8]), .b(b[11:8]), .cin(out[1]), .cout(out[2]), .sum(sum[11:8]));
    bcd_fadd_diy bcd_fadd3 (.a(a[15:12]), .b(b[15:12]), .cin(out[2]), .cout(cout), .sum(sum[15:12]));
`else
    bcd_fadd bcd_fadd0 (.a(a[3:0]), .b(b[3:0]), .cin(cin), .cout(out[0]), .sum(sum[3:0]));
    bcd_fadd bcd_fadd1 (.a(a[7:4]), .b(b[7:4]), .cin(out[0]), .cout(out[1]), .sum(sum[7:4]));
    bcd_fadd bcd_fadd2 (.a(a[11:8]), .b(b[11:8]), .cin(out[1]), .cout(out[2]), .sum(sum[11:8]));
    bcd_fadd bcd_fadd3 (.a(a[15:12]), .b(b[15:12]), .cin(out[2]), .cout(cout), .sum(sum[15:12]));
`endif
endmodule

module bcd_fadd_diy ( 
    input [3:0] a, b,
    input cin,
    output cout,
    output [3:0] sum );
    
    wire cout0, cout1;
    wire [3:0] sum0, sum1;
    localparam ANS_SEL = 0;
    assign {cout, sum} = ANS_SEL ? {cout1, sum1} : {cout0, sum0};
    // method1
    wire [5:0] sum_temp = cin + a + b;
    assign cout0 = sum_temp > 'd9;
    assign sum0 = cout ? sum_temp - 'd10 : sum_temp;
    // method2
    always @ (*) begin
        case({cin, b, a})
        'h000: {cout1, sum1} = 'h00;
        'h001: {cout1, sum1} = 'h01;
        'h002: {cout1, sum1} = 'h02;
        'h003: {cout1, sum1} = 'h03;
        'h004: {cout1, sum1} = 'h04;
        'h005: {cout1, sum1} = 'h05;
        'h006: {cout1, sum1} = 'h06;
        'h007: {cout1, sum1} = 'h07;
        'h008: {cout1, sum1} = 'h08;
        'h009: {cout1, sum1} = 'h09;
        'h00A: {cout1, sum1} = 'h10;
        'h00B: {cout1, sum1} = 'h11;
        'h00C: {cout1, sum1} = 'h12;
        'h00D: {cout1, sum1} = 'h13;
        'h00E: {cout1, sum1} = 'h14;
        'h00F: {cout1, sum1} = 'h15;
        'h010: {cout1, sum1} = 'h01;
        'h011: {cout1, sum1} = 'h02;
        'h012: {cout1, sum1} = 'h03;
        'h013: {cout1, sum1} = 'h04;
        'h014: {cout1, sum1} = 'h05;
        'h015: {cout1, sum1} = 'h06;
        'h016: {cout1, sum1} = 'h07;
        'h017: {cout1, sum1} = 'h08;
        'h018: {cout1, sum1} = 'h09;
        'h019: {cout1, sum1} = 'h10;
        'h01A: {cout1, sum1} = 'h11;
        'h01B: {cout1, sum1} = 'h12;
        'h01C: {cout1, sum1} = 'h13;
        'h01D: {cout1, sum1} = 'h14;
        'h01E: {cout1, sum1} = 'h15;
        'h01F: {cout1, sum1} = 'h16;
        'h020: {cout1, sum1} = 'h02;
        'h021: {cout1, sum1} = 'h03;
        'h022: {cout1, sum1} = 'h04;
        'h023: {cout1, sum1} = 'h05;
        'h024: {cout1, sum1} = 'h06;
        'h025: {cout1, sum1} = 'h07;
        'h026: {cout1, sum1} = 'h08;
        'h027: {cout1, sum1} = 'h09;
        'h028: {cout1, sum1} = 'h10;
        'h029: {cout1, sum1} = 'h11;
        'h02A: {cout1, sum1} = 'h12;
        'h02B: {cout1, sum1} = 'h13;
        'h02C: {cout1, sum1} = 'h14;
        'h02D: {cout1, sum1} = 'h15;
        'h02E: {cout1, sum1} = 'h16;
        'h02F: {cout1, sum1} = 'h17;
        'h030: {cout1, sum1} = 'h03;
        'h031: {cout1, sum1} = 'h04;
        'h032: {cout1, sum1} = 'h05;
        'h033: {cout1, sum1} = 'h06;
        'h034: {cout1, sum1} = 'h07;
        'h035: {cout1, sum1} = 'h08;
        'h036: {cout1, sum1} = 'h09;
        'h037: {cout1, sum1} = 'h10;
        'h038: {cout1, sum1} = 'h11;
        'h039: {cout1, sum1} = 'h12;
        'h03A: {cout1, sum1} = 'h13;
        'h03B: {cout1, sum1} = 'h14;
        'h03C: {cout1, sum1} = 'h15;
        'h03D: {cout1, sum1} = 'h16;
        'h03E: {cout1, sum1} = 'h17;
        'h03F: {cout1, sum1} = 'h18;
        'h040: {cout1, sum1} = 'h04;
        'h041: {cout1, sum1} = 'h05;
        'h042: {cout1, sum1} = 'h06;
        'h043: {cout1, sum1} = 'h07;
        'h044: {cout1, sum1} = 'h08;
        'h045: {cout1, sum1} = 'h09;
        'h046: {cout1, sum1} = 'h10;
        'h047: {cout1, sum1} = 'h11;
        'h048: {cout1, sum1} = 'h12;
        'h049: {cout1, sum1} = 'h13;
        'h04A: {cout1, sum1} = 'h14;
        'h04B: {cout1, sum1} = 'h15;
        'h04C: {cout1, sum1} = 'h16;
        'h04D: {cout1, sum1} = 'h17;
        'h04E: {cout1, sum1} = 'h18;
        'h04F: {cout1, sum1} = 'h19;
        'h050: {cout1, sum1} = 'h05;
        'h051: {cout1, sum1} = 'h06;
        'h052: {cout1, sum1} = 'h07;
        'h053: {cout1, sum1} = 'h08;
        'h054: {cout1, sum1} = 'h09;
        'h055: {cout1, sum1} = 'h10;
        'h056: {cout1, sum1} = 'h11;
        'h057: {cout1, sum1} = 'h12;
        'h058: {cout1, sum1} = 'h13;
        'h059: {cout1, sum1} = 'h14;
        'h05A: {cout1, sum1} = 'h15;
        'h05B: {cout1, sum1} = 'h16;
        'h05C: {cout1, sum1} = 'h17;
        'h05D: {cout1, sum1} = 'h18;
        'h05E: {cout1, sum1} = 'h19;
        'h05F: {cout1, sum1} = 'h10;
        'h060: {cout1, sum1} = 'h06;
        'h061: {cout1, sum1} = 'h07;
        'h062: {cout1, sum1} = 'h08;
        'h063: {cout1, sum1} = 'h09;
        'h064: {cout1, sum1} = 'h10;
        'h065: {cout1, sum1} = 'h11;
        'h066: {cout1, sum1} = 'h12;
        'h067: {cout1, sum1} = 'h13;
        'h068: {cout1, sum1} = 'h14;
        'h069: {cout1, sum1} = 'h15;
        'h06A: {cout1, sum1} = 'h16;
        'h06B: {cout1, sum1} = 'h17;
        'h06C: {cout1, sum1} = 'h18;
        'h06D: {cout1, sum1} = 'h19;
        'h06E: {cout1, sum1} = 'h10;
        'h06F: {cout1, sum1} = 'h11;
        'h070: {cout1, sum1} = 'h07;
        'h071: {cout1, sum1} = 'h08;
        'h072: {cout1, sum1} = 'h09;
        'h073: {cout1, sum1} = 'h10;
        'h074: {cout1, sum1} = 'h11;
        'h075: {cout1, sum1} = 'h12;
        'h076: {cout1, sum1} = 'h13;
        'h077: {cout1, sum1} = 'h14;
        'h078: {cout1, sum1} = 'h15;
        'h079: {cout1, sum1} = 'h16;
        'h07A: {cout1, sum1} = 'h17;
        'h07B: {cout1, sum1} = 'h18;
        'h07C: {cout1, sum1} = 'h19;
        'h07D: {cout1, sum1} = 'h10;
        'h07E: {cout1, sum1} = 'h11;
        'h07F: {cout1, sum1} = 'h12;
        'h080: {cout1, sum1} = 'h08;
        'h081: {cout1, sum1} = 'h09;
        'h082: {cout1, sum1} = 'h10;
        'h083: {cout1, sum1} = 'h11;
        'h084: {cout1, sum1} = 'h12;
        'h085: {cout1, sum1} = 'h13;
        'h086: {cout1, sum1} = 'h14;
        'h087: {cout1, sum1} = 'h15;
        'h088: {cout1, sum1} = 'h16;
        'h089: {cout1, sum1} = 'h17;
        'h08A: {cout1, sum1} = 'h18;
        'h08B: {cout1, sum1} = 'h19;
        'h08C: {cout1, sum1} = 'h10;
        'h08D: {cout1, sum1} = 'h11;
        'h08E: {cout1, sum1} = 'h12;
        'h08F: {cout1, sum1} = 'h13;
        'h090: {cout1, sum1} = 'h09;
        'h091: {cout1, sum1} = 'h10;
        'h092: {cout1, sum1} = 'h11;
        'h093: {cout1, sum1} = 'h12;
        'h094: {cout1, sum1} = 'h13;
        'h095: {cout1, sum1} = 'h14;
        'h096: {cout1, sum1} = 'h15;
        'h097: {cout1, sum1} = 'h16;
        'h098: {cout1, sum1} = 'h17;
        'h099: {cout1, sum1} = 'h18;
        'h09A: {cout1, sum1} = 'h19;
        'h09B: {cout1, sum1} = 'h10;
        'h09C: {cout1, sum1} = 'h11;
        'h09D: {cout1, sum1} = 'h12;
        'h09E: {cout1, sum1} = 'h13;
        'h09F: {cout1, sum1} = 'h14;
        'h0A0: {cout1, sum1} = 'h10;
        'h0A1: {cout1, sum1} = 'h11;
        'h0A2: {cout1, sum1} = 'h12;
        'h0A3: {cout1, sum1} = 'h13;
        'h0A4: {cout1, sum1} = 'h14;
        'h0A5: {cout1, sum1} = 'h15;
        'h0A6: {cout1, sum1} = 'h16;
        'h0A7: {cout1, sum1} = 'h17;
        'h0A8: {cout1, sum1} = 'h18;
        'h0A9: {cout1, sum1} = 'h19;
        'h0AA: {cout1, sum1} = 'h10;
        'h0AB: {cout1, sum1} = 'h11;
        'h0AC: {cout1, sum1} = 'h12;
        'h0AD: {cout1, sum1} = 'h13;
        'h0AE: {cout1, sum1} = 'h14;
        'h0AF: {cout1, sum1} = 'h15;
        'h0B0: {cout1, sum1} = 'h11;
        'h0B1: {cout1, sum1} = 'h12;
        'h0B2: {cout1, sum1} = 'h13;
        'h0B3: {cout1, sum1} = 'h14;
        'h0B4: {cout1, sum1} = 'h15;
        'h0B5: {cout1, sum1} = 'h16;
        'h0B6: {cout1, sum1} = 'h17;
        'h0B7: {cout1, sum1} = 'h18;
        'h0B8: {cout1, sum1} = 'h19;
        'h0B9: {cout1, sum1} = 'h10;
        'h0BA: {cout1, sum1} = 'h11;
        'h0BB: {cout1, sum1} = 'h12;
        'h0BC: {cout1, sum1} = 'h13;
        'h0BD: {cout1, sum1} = 'h14;
        'h0BE: {cout1, sum1} = 'h15;
        'h0BF: {cout1, sum1} = 'h16;
        'h0C0: {cout1, sum1} = 'h12;
        'h0C1: {cout1, sum1} = 'h13;
        'h0C2: {cout1, sum1} = 'h14;
        'h0C3: {cout1, sum1} = 'h15;
        'h0C4: {cout1, sum1} = 'h16;
        'h0C5: {cout1, sum1} = 'h17;
        'h0C6: {cout1, sum1} = 'h18;
        'h0C7: {cout1, sum1} = 'h19;
        'h0C8: {cout1, sum1} = 'h10;
        'h0C9: {cout1, sum1} = 'h11;
        'h0CA: {cout1, sum1} = 'h12;
        'h0CB: {cout1, sum1} = 'h13;
        'h0CC: {cout1, sum1} = 'h14;
        'h0CD: {cout1, sum1} = 'h15;
        'h0CE: {cout1, sum1} = 'h16;
        'h0CF: {cout1, sum1} = 'h17;
        'h0D0: {cout1, sum1} = 'h13;
        'h0D1: {cout1, sum1} = 'h14;
        'h0D2: {cout1, sum1} = 'h15;
        'h0D3: {cout1, sum1} = 'h16;
        'h0D4: {cout1, sum1} = 'h17;
        'h0D5: {cout1, sum1} = 'h18;
        'h0D6: {cout1, sum1} = 'h19;
        'h0D7: {cout1, sum1} = 'h10;
        'h0D8: {cout1, sum1} = 'h11;
        'h0D9: {cout1, sum1} = 'h12;
        'h0DA: {cout1, sum1} = 'h13;
        'h0DB: {cout1, sum1} = 'h14;
        'h0DC: {cout1, sum1} = 'h15;
        'h0DD: {cout1, sum1} = 'h16;
        'h0DE: {cout1, sum1} = 'h17;
        'h0DF: {cout1, sum1} = 'h18;
        'h0E0: {cout1, sum1} = 'h14;
        'h0E1: {cout1, sum1} = 'h15;
        'h0E2: {cout1, sum1} = 'h16;
        'h0E3: {cout1, sum1} = 'h17;
        'h0E4: {cout1, sum1} = 'h18;
        'h0E5: {cout1, sum1} = 'h19;
        'h0E6: {cout1, sum1} = 'h10;
        'h0E7: {cout1, sum1} = 'h11;
        'h0E8: {cout1, sum1} = 'h12;
        'h0E9: {cout1, sum1} = 'h13;
        'h0EA: {cout1, sum1} = 'h14;
        'h0EB: {cout1, sum1} = 'h15;
        'h0EC: {cout1, sum1} = 'h16;
        'h0ED: {cout1, sum1} = 'h17;
        'h0EE: {cout1, sum1} = 'h18;
        'h0EF: {cout1, sum1} = 'h19;
        'h0F0: {cout1, sum1} = 'h15;
        'h0F1: {cout1, sum1} = 'h16;
        'h0F2: {cout1, sum1} = 'h17;
        'h0F3: {cout1, sum1} = 'h18;
        'h0F4: {cout1, sum1} = 'h19;
        'h0F5: {cout1, sum1} = 'h10;
        'h0F6: {cout1, sum1} = 'h11;
        'h0F7: {cout1, sum1} = 'h12;
        'h0F8: {cout1, sum1} = 'h13;
        'h0F9: {cout1, sum1} = 'h14;
        'h0FA: {cout1, sum1} = 'h15;
        'h0FB: {cout1, sum1} = 'h16;
        'h0FC: {cout1, sum1} = 'h17;
        'h0FD: {cout1, sum1} = 'h18;
        'h0FE: {cout1, sum1} = 'h19;
        'h0FF: {cout1, sum1} = 'h10;
        'h100: {cout1, sum1} = 'h01;
        'h101: {cout1, sum1} = 'h02;
        'h102: {cout1, sum1} = 'h03;
        'h103: {cout1, sum1} = 'h04;
        'h104: {cout1, sum1} = 'h05;
        'h105: {cout1, sum1} = 'h06;
        'h106: {cout1, sum1} = 'h07;
        'h107: {cout1, sum1} = 'h08;
        'h108: {cout1, sum1} = 'h09;
        'h109: {cout1, sum1} = 'h10;
        'h10A: {cout1, sum1} = 'h11;
        'h10B: {cout1, sum1} = 'h12;
        'h10C: {cout1, sum1} = 'h13;
        'h10D: {cout1, sum1} = 'h14;
        'h10E: {cout1, sum1} = 'h15;
        'h10F: {cout1, sum1} = 'h16;
        'h110: {cout1, sum1} = 'h02;
        'h111: {cout1, sum1} = 'h03;
        'h112: {cout1, sum1} = 'h04;
        'h113: {cout1, sum1} = 'h05;
        'h114: {cout1, sum1} = 'h06;
        'h115: {cout1, sum1} = 'h07;
        'h116: {cout1, sum1} = 'h08;
        'h117: {cout1, sum1} = 'h09;
        'h118: {cout1, sum1} = 'h10;
        'h119: {cout1, sum1} = 'h11;
        'h11A: {cout1, sum1} = 'h12;
        'h11B: {cout1, sum1} = 'h13;
        'h11C: {cout1, sum1} = 'h14;
        'h11D: {cout1, sum1} = 'h15;
        'h11E: {cout1, sum1} = 'h16;
        'h11F: {cout1, sum1} = 'h17;
        'h120: {cout1, sum1} = 'h03;
        'h121: {cout1, sum1} = 'h04;
        'h122: {cout1, sum1} = 'h05;
        'h123: {cout1, sum1} = 'h06;
        'h124: {cout1, sum1} = 'h07;
        'h125: {cout1, sum1} = 'h08;
        'h126: {cout1, sum1} = 'h09;
        'h127: {cout1, sum1} = 'h10;
        'h128: {cout1, sum1} = 'h11;
        'h129: {cout1, sum1} = 'h12;
        'h12A: {cout1, sum1} = 'h13;
        'h12B: {cout1, sum1} = 'h14;
        'h12C: {cout1, sum1} = 'h15;
        'h12D: {cout1, sum1} = 'h16;
        'h12E: {cout1, sum1} = 'h17;
        'h12F: {cout1, sum1} = 'h18;
        'h130: {cout1, sum1} = 'h04;
        'h131: {cout1, sum1} = 'h05;
        'h132: {cout1, sum1} = 'h06;
        'h133: {cout1, sum1} = 'h07;
        'h134: {cout1, sum1} = 'h08;
        'h135: {cout1, sum1} = 'h09;
        'h136: {cout1, sum1} = 'h10;
        'h137: {cout1, sum1} = 'h11;
        'h138: {cout1, sum1} = 'h12;
        'h139: {cout1, sum1} = 'h13;
        'h13A: {cout1, sum1} = 'h14;
        'h13B: {cout1, sum1} = 'h15;
        'h13C: {cout1, sum1} = 'h16;
        'h13D: {cout1, sum1} = 'h17;
        'h13E: {cout1, sum1} = 'h18;
        'h13F: {cout1, sum1} = 'h19;
        'h140: {cout1, sum1} = 'h05;
        'h141: {cout1, sum1} = 'h06;
        'h142: {cout1, sum1} = 'h07;
        'h143: {cout1, sum1} = 'h08;
        'h144: {cout1, sum1} = 'h09;
        'h145: {cout1, sum1} = 'h10;
        'h146: {cout1, sum1} = 'h11;
        'h147: {cout1, sum1} = 'h12;
        'h148: {cout1, sum1} = 'h13;
        'h149: {cout1, sum1} = 'h14;
        'h14A: {cout1, sum1} = 'h15;
        'h14B: {cout1, sum1} = 'h16;
        'h14C: {cout1, sum1} = 'h17;
        'h14D: {cout1, sum1} = 'h18;
        'h14E: {cout1, sum1} = 'h19;
        'h14F: {cout1, sum1} = 'h10;
        'h150: {cout1, sum1} = 'h06;
        'h151: {cout1, sum1} = 'h07;
        'h152: {cout1, sum1} = 'h08;
        'h153: {cout1, sum1} = 'h09;
        'h154: {cout1, sum1} = 'h10;
        'h155: {cout1, sum1} = 'h11;
        'h156: {cout1, sum1} = 'h12;
        'h157: {cout1, sum1} = 'h13;
        'h158: {cout1, sum1} = 'h14;
        'h159: {cout1, sum1} = 'h15;
        'h15A: {cout1, sum1} = 'h16;
        'h15B: {cout1, sum1} = 'h17;
        'h15C: {cout1, sum1} = 'h18;
        'h15D: {cout1, sum1} = 'h19;
        'h15E: {cout1, sum1} = 'h10;
        'h15F: {cout1, sum1} = 'h11;
        'h160: {cout1, sum1} = 'h07;
        'h161: {cout1, sum1} = 'h08;
        'h162: {cout1, sum1} = 'h09;
        'h163: {cout1, sum1} = 'h10;
        'h164: {cout1, sum1} = 'h11;
        'h165: {cout1, sum1} = 'h12;
        'h166: {cout1, sum1} = 'h13;
        'h167: {cout1, sum1} = 'h14;
        'h168: {cout1, sum1} = 'h15;
        'h169: {cout1, sum1} = 'h16;
        'h16A: {cout1, sum1} = 'h17;
        'h16B: {cout1, sum1} = 'h18;
        'h16C: {cout1, sum1} = 'h19;
        'h16D: {cout1, sum1} = 'h10;
        'h16E: {cout1, sum1} = 'h11;
        'h16F: {cout1, sum1} = 'h12;
        'h170: {cout1, sum1} = 'h08;
        'h171: {cout1, sum1} = 'h09;
        'h172: {cout1, sum1} = 'h10;
        'h173: {cout1, sum1} = 'h11;
        'h174: {cout1, sum1} = 'h12;
        'h175: {cout1, sum1} = 'h13;
        'h176: {cout1, sum1} = 'h14;
        'h177: {cout1, sum1} = 'h15;
        'h178: {cout1, sum1} = 'h16;
        'h179: {cout1, sum1} = 'h17;
        'h17A: {cout1, sum1} = 'h18;
        'h17B: {cout1, sum1} = 'h19;
        'h17C: {cout1, sum1} = 'h10;
        'h17D: {cout1, sum1} = 'h11;
        'h17E: {cout1, sum1} = 'h12;
        'h17F: {cout1, sum1} = 'h13;
        'h180: {cout1, sum1} = 'h09;
        'h181: {cout1, sum1} = 'h10;
        'h182: {cout1, sum1} = 'h11;
        'h183: {cout1, sum1} = 'h12;
        'h184: {cout1, sum1} = 'h13;
        'h185: {cout1, sum1} = 'h14;
        'h186: {cout1, sum1} = 'h15;
        'h187: {cout1, sum1} = 'h16;
        'h188: {cout1, sum1} = 'h17;
        'h189: {cout1, sum1} = 'h18;
        'h18A: {cout1, sum1} = 'h19;
        'h18B: {cout1, sum1} = 'h10;
        'h18C: {cout1, sum1} = 'h11;
        'h18D: {cout1, sum1} = 'h12;
        'h18E: {cout1, sum1} = 'h13;
        'h18F: {cout1, sum1} = 'h14;
        'h190: {cout1, sum1} = 'h10;
        'h191: {cout1, sum1} = 'h11;
        'h192: {cout1, sum1} = 'h12;
        'h193: {cout1, sum1} = 'h13;
        'h194: {cout1, sum1} = 'h14;
        'h195: {cout1, sum1} = 'h15;
        'h196: {cout1, sum1} = 'h16;
        'h197: {cout1, sum1} = 'h17;
        'h198: {cout1, sum1} = 'h18;
        'h199: {cout1, sum1} = 'h19;
        'h19A: {cout1, sum1} = 'h10;
        'h19B: {cout1, sum1} = 'h11;
        'h19C: {cout1, sum1} = 'h12;
        'h19D: {cout1, sum1} = 'h13;
        'h19E: {cout1, sum1} = 'h14;
        'h19F: {cout1, sum1} = 'h15;
        'h1A0: {cout1, sum1} = 'h11;
        'h1A1: {cout1, sum1} = 'h12;
        'h1A2: {cout1, sum1} = 'h13;
        'h1A3: {cout1, sum1} = 'h14;
        'h1A4: {cout1, sum1} = 'h15;
        'h1A5: {cout1, sum1} = 'h16;
        'h1A6: {cout1, sum1} = 'h17;
        'h1A7: {cout1, sum1} = 'h18;
        'h1A8: {cout1, sum1} = 'h19;
        'h1A9: {cout1, sum1} = 'h10;
        'h1AA: {cout1, sum1} = 'h11;
        'h1AB: {cout1, sum1} = 'h12;
        'h1AC: {cout1, sum1} = 'h13;
        'h1AD: {cout1, sum1} = 'h14;
        'h1AE: {cout1, sum1} = 'h15;
        'h1AF: {cout1, sum1} = 'h16;
        'h1B0: {cout1, sum1} = 'h12;
        'h1B1: {cout1, sum1} = 'h13;
        'h1B2: {cout1, sum1} = 'h14;
        'h1B3: {cout1, sum1} = 'h15;
        'h1B4: {cout1, sum1} = 'h16;
        'h1B5: {cout1, sum1} = 'h17;
        'h1B6: {cout1, sum1} = 'h18;
        'h1B7: {cout1, sum1} = 'h19;
        'h1B8: {cout1, sum1} = 'h10;
        'h1B9: {cout1, sum1} = 'h11;
        'h1BA: {cout1, sum1} = 'h12;
        'h1BB: {cout1, sum1} = 'h13;
        'h1BC: {cout1, sum1} = 'h14;
        'h1BD: {cout1, sum1} = 'h15;
        'h1BE: {cout1, sum1} = 'h16;
        'h1BF: {cout1, sum1} = 'h17;
        'h1C0: {cout1, sum1} = 'h13;
        'h1C1: {cout1, sum1} = 'h14;
        'h1C2: {cout1, sum1} = 'h15;
        'h1C3: {cout1, sum1} = 'h16;
        'h1C4: {cout1, sum1} = 'h17;
        'h1C5: {cout1, sum1} = 'h18;
        'h1C6: {cout1, sum1} = 'h19;
        'h1C7: {cout1, sum1} = 'h10;
        'h1C8: {cout1, sum1} = 'h11;
        'h1C9: {cout1, sum1} = 'h12;
        'h1CA: {cout1, sum1} = 'h13;
        'h1CB: {cout1, sum1} = 'h14;
        'h1CC: {cout1, sum1} = 'h15;
        'h1CD: {cout1, sum1} = 'h16;
        'h1CE: {cout1, sum1} = 'h17;
        'h1CF: {cout1, sum1} = 'h18;
        'h1D0: {cout1, sum1} = 'h14;
        'h1D1: {cout1, sum1} = 'h15;
        'h1D2: {cout1, sum1} = 'h16;
        'h1D3: {cout1, sum1} = 'h17;
        'h1D4: {cout1, sum1} = 'h18;
        'h1D5: {cout1, sum1} = 'h19;
        'h1D6: {cout1, sum1} = 'h10;
        'h1D7: {cout1, sum1} = 'h11;
        'h1D8: {cout1, sum1} = 'h12;
        'h1D9: {cout1, sum1} = 'h13;
        'h1DA: {cout1, sum1} = 'h14;
        'h1DB: {cout1, sum1} = 'h15;
        'h1DC: {cout1, sum1} = 'h16;
        'h1DD: {cout1, sum1} = 'h17;
        'h1DE: {cout1, sum1} = 'h18;
        'h1DF: {cout1, sum1} = 'h19;
        'h1E0: {cout1, sum1} = 'h15;
        'h1E1: {cout1, sum1} = 'h16;
        'h1E2: {cout1, sum1} = 'h17;
        'h1E3: {cout1, sum1} = 'h18;
        'h1E4: {cout1, sum1} = 'h19;
        'h1E5: {cout1, sum1} = 'h10;
        'h1E6: {cout1, sum1} = 'h11;
        'h1E7: {cout1, sum1} = 'h12;
        'h1E8: {cout1, sum1} = 'h13;
        'h1E9: {cout1, sum1} = 'h14;
        'h1EA: {cout1, sum1} = 'h15;
        'h1EB: {cout1, sum1} = 'h16;
        'h1EC: {cout1, sum1} = 'h17;
        'h1ED: {cout1, sum1} = 'h18;
        'h1EE: {cout1, sum1} = 'h19;
        'h1EF: {cout1, sum1} = 'h10;
        'h1F0: {cout1, sum1} = 'h16;
        'h1F1: {cout1, sum1} = 'h17;
        'h1F2: {cout1, sum1} = 'h18;
        'h1F3: {cout1, sum1} = 'h19;
        'h1F4: {cout1, sum1} = 'h10;
        'h1F5: {cout1, sum1} = 'h11;
        'h1F6: {cout1, sum1} = 'h12;
        'h1F7: {cout1, sum1} = 'h13;
        'h1F8: {cout1, sum1} = 'h14;
        'h1F9: {cout1, sum1} = 'h15;
        'h1FA: {cout1, sum1} = 'h16;
        'h1FB: {cout1, sum1} = 'h17;
        'h1FC: {cout1, sum1} = 'h18;
        'h1FD: {cout1, sum1} = 'h19;
        'h1FE: {cout1, sum1} = 'h10;
        'h1FF: {cout1, sum1} = 'h11;
        endcase
    end
endmodule
