module top_module_p165 ();
endmodule
