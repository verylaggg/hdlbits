module top_module_p91 ();
endmodule
