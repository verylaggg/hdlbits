module top_module_p60 ();
endmodule
