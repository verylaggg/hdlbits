module top_module_p62 ();
endmodule
