module top_module_p47 ();
endmodule
